
module tarea1 (
	clk_clk);	

	input		clk_clk;
endmodule
